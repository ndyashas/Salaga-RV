`ifndef CORE_VARIANT

`define CORE_VARIANT eka


`endif
