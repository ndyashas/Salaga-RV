`ifndef CORE_VARIANT

`define CORE_VARIANT eka

/*
 * Each of l1 data and instruction caches
 * are of size 16Kbytes
 */
`define CACHE_ADDRESS_SIZE 14

`endif
